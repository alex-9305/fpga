`include "windows_fsm.v"
`timescale 1us/1ns

module windows_fsm_tb


endmodule