module i2c_master
    (

    );



endmodule